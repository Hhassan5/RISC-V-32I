`timescale 1ns / 1ps



module InstMem#(n=32)(
input [5:0] addr,
output [n-1:0] data_out
);
    reg [n-1:0] mem [0:63];
    
    assign data_out = mem[addr];
    

initial begin
mem[0]=32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0) 
mem[1]=32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0) 
mem[2]=32'b01000000001000001000000110110011 ; //sub x3, x1, x2 
mem[3]=32'b00000000001000001000001000110011 ; //add x4, x1, x2 
mem[4]=32'b00000000001000001000010001100011 ; //beq x1, x2, 8  
mem[5]=32'b01000000001000001000000110110011 ; //sub x3, x1, x
mem[6]=32'b00000000010000001111001010110011 ; //and x5, x1, x4 
mem[7]=32'b00000000001000001011010000110011;//sltu x8, x1, x2
mem[8]=32'b00000000001000001010010010110011;//slt x9, x1, x2
mem[9]=32'b00000000001000001101010100110011;//srl x10, x1, x2
mem[10]=32'b00000000001000001001010110110011;//sll x11, x1, x2
mem[11]=32'b01000000000100010000011000110011;//sub x12, x2, x1

mem[12]=32'b00000000001100001111011010010011;//andi x13, x1, 3 
mem[13]=32'b00000000001100001110011100010011;//ori x14, x1, 3
mem[14]=32'b00000000001100001100011110010011;//xori x15, x1, 3 
mem[15]=32'b00000000001100001011100000010011;//sltiu x16, x1, 3 
mem[16]=32'b11111111110100001010100010010011;//slti x17, x1, -3
mem[17]=32'b00000000001100001000100100010011;//addi x18, x1, 3

mem[18]=32'b00000000000000001010100110010111;//auipc x19,10 
mem[19]=32'b00000000000000001010101000110111;//lui x20,10 


//mem[20]=32'b00000000000000001000101101100111;//jalr x22, 0(x1) 
//mem[21]=32'b00000000010000000000101111101111;//jal x23, 4 
mem[22]=32'b00000000001000001010000000100011;//sw x2, 0(x1) 

//Branch
mem[23]=32'b00000000001000001111001001100011;//bgeu x1, x2, 4
mem[24]=32'b00000000001000001110010001100011;//bltu x1, x2, 8 
mem[25]=32'b00000000001000001101001001100011;//bge x1, x2, 4 
mem[26]=32'b00000000001000001100010001100011;//blt x1, x2, 8 
mem[27]=32'b00000000001000001001001001100011;//bne x1, x2, 4 
mem[28]=32'b00000000010100010000011001100011;//beq x1, x2, 8 

//mem[40]=32'b00000000010100001001000000100011; //sh x17, 0(x1) 
//mem[41]=32'b00000000010100001000000000100011; //sb x12, 0(x2) 
//mem[42]=32'b00000000100000000101000110000011;//lhu x13, 0(x1) 
//mem[43]=32'b00000000100000000100000110000011;//lbu x14, 0(x2)
//mem[44]=32'b00000000100000000000000110000011;//lb x15, 0(x1) 
//mem[45]=32'b00000000100000000001000110000011;// lh x16, 0(x2)     
   
    end
    
endmodule

